//==============================================================================
//  Filename    : bench_riscv
//  Description : General test bench for the RISC-V processor
//==============================================================================

module bench_riscv();

timeunit      1ns;
timeprecision 1ns;

// Simulation parameters
localparam  MEM_SIZE   = 4095, 
            PROG_SIZE  = 683,
            CLK_PERIOD = 20, 
            NB_TESTS   = 292/*25*/;

logic [31:0]  insn_buff[PROG_SIZE:0];                       // Buffer to read

int clock_number;                                           // Number of clock cycles since the reset
int passed_test = 0;                                        // Number of passed tests
int done_test = 0;                                          // Number of done tests
int value_ok = 0;                                           // Inidicate if the value read is the expected one

typedef struct {
    string name;
    int clk;
    logic [32:0] address;
    int size;
    logic [31:0] value;
} tests;

// Test cases : See asm_bench_global.xlsx for more details
//                         name,                    clk,  address, size, value
/*tests test[NB_TESTS] = '{'{"ADD sans débordement ", 26,   22     ,  8,   32'h0000001E},
                         '{"ADD avec débordement ", 30,   4      , 32,   32'h0F0F070D},
                         '{"AND                  ", 51,   4      , 32,   32'h0F0F070E},
                         '{"SLL                  ", 72,   16     , 16,   32'h00000000},
                         '{"SRL                  ", 93,   16     , 16,   32'h00000001},
                         '{"OR                   ", 114,  4      , 32,   32'hFFFFFFFF},
                         '{"XOR                  ", 135,  4      , 32,   32'hF0F0F8F1},
                         '{"SLTU true            ", 157,  22     , 8,    32'h00000001},
                         '{"SLTU false           ", 162,  16     , 16,   32'h00000000},
                         '{"SLT true             ", 184,  22     , 8,    32'h00000001},
                         '{"SLT false            ", 189,  16     , 16,   32'h00000000},
                         '{"SRA                  ", 210,  16     , 16,   32'h00000001},
                         '{"SUB sans débordement ", 231,  22     , 8,    32'h00000001},
                         '{"SUB avec débordement ", 235,  16     , 16,   32'hFFFF0011},
                         '{"SLLI avec débordement", 255,  16     , 16,   32'h0000FFC0},
                         '{"SLLI sans débordement", 258,  22     , 8,    32'h000000C0},
                         '{"SRLI sans débordement", 278,  31     , 16,   32'h00007F87},
                         '{"SRLI avec débordement", 281,  22     , 8,    32'h00000010},
                         '{"ORI                  ", 303,  4      , 32,   32'h0000070F},
                         '{"ORI  avec dépendance ", 304,  8      , 32,   32'hFFFFFFFF},
                         '{"XORI                 ", 326,  4      , 32,   32'hF0F0F8F1},
                         '{"SLTIU true           ", 350,  22     , 8,    32'h00000001},
                         '{"SLTIU false          ", 354,  16     , 16,   32'h00000000},
                         '{"SLTI true            ", 375,  22     , 16,   32'h00000001},
                         '{"SLTI false           ", 379,  16     , 16,   32'h00000000}/*,
                         TODO : tests sur les branchements*/
                    //    };

tests test[NB_TESTS] = '{
'{"PC = 4 : SW", 1, 48, 32, 32'h00000000},              // 00004 sw     fp,48(sp)
'{"PC = 40 : SB", 10, 2755, 8, 32'h0000000e},           // 00040 sb     a5,-17(fp)
'{"PC = 48 : SB", 12, 2747, 8, 32'h0000000f},           // 00048 sb     a5,-25(fp)
'{"PC = 56 : SB", 14, 2746, 8, 32'h00000001},           // 00056 sb     a5,-26(fp)
'{"PC = 64 : SH", 16, 2744, 16, 32'hfffffffe},          // 00064 sh     a5,-28(fp)
'{"PC = 72 : SH", 18, 2742, 16, 32'h0000000f},          // 00072 sh     a5,-30(fp)
'{"PC = 76 : SH", 19, 2740, 16, 32'h00000000},          // 00076 sh     zero,-32(fp)
'{"PC = 84 : SW", 21, 2736, 32, 32'hfffffffe},          // 00084 sw     a5,-36(fp)
'{"PC = 96 : SW", 24, 2732, 32, 32'h0f0f070f},          // 00096 sw     a5,-40(fp)
'{"PC = 100 : SW", 25, 2728, 32, 32'h00000000},         // 00100 sw     zero,-44(fp)
'{"PC = 128 : SB", 32, 2746, 8, 32'h0000001e},          // 00128 sb     a5,-26(fp)
'{"PC = 144 : SW", 36, 2728, 32, 32'h0f0f070d},         // 00144 sw     a5,-44(fp)
'{"PC = 152 : SB", 38, 2755, 8, 32'h0000000e},          // 00152 sb     a5,-17(fp)
'{"PC = 160 : SB", 40, 2747, 8, 32'h0000000f},          // 00160 sb     a5,-25(fp)
'{"PC = 168 : SB", 42, 2746, 8, 32'h00000001},          // 00168 sb     a5,-26(fp)
'{"PC = 176 : SH", 44, 2744, 16, 32'hfffffffe},         // 00176 sh     a5,-28(fp)
'{"PC = 184 : SH", 46, 2742, 16, 32'h0000000f},         // 00184 sh     a5,-30(fp)
'{"PC = 188 : SH", 47, 2740, 16, 32'h00000000},         // 00188 sh     zero,-32(fp)
'{"PC = 196 : SW", 49, 2736, 32, 32'hfffffffe},         // 00196 sw     a5,-36(fp)
'{"PC = 208 : SW", 52, 2732, 32, 32'h0f0f070f},         // 00208 sw     a5,-40(fp)
'{"PC = 212 : SW", 53, 2728, 32, 32'h00000000},         // 00212 sw     zero,-44(fp)
'{"PC = 228 : SW", 57, 2728, 32, 32'h0f0f070e},         // 00228 sw     a5,-44(fp)
'{"PC = 236 : SB", 59, 2755, 8, 32'h0000000e},          // 00236 sb     a5,-17(fp)
'{"PC = 244 : SB", 61, 2747, 8, 32'h0000000f},          // 00244 sb     a5,-25(fp)
'{"PC = 252 : SB", 63, 2746, 8, 32'h00000001},          // 00252 sb     a5,-26(fp)
'{"PC = 260 : SH", 65, 2744, 16, 32'hfffffffe},         // 00260 sh     a5,-28(fp)
'{"PC = 268 : SH", 67, 2742, 16, 32'h0000000f},         // 00268 sh     a5,-30(fp)
'{"PC = 272 : SH", 68, 2740, 16, 32'h00000000},         // 00272 sh     zero,-32(fp)
'{"PC = 280 : SW", 70, 2736, 32, 32'hfffffffe},         // 00280 sw     a5,-36(fp)
'{"PC = 292 : SW", 73, 2732, 32, 32'h0f0f070f},         // 00292 sw     a5,-40(fp)
'{"PC = 296 : SW", 74, 2728, 32, 32'h00000000},         // 00296 sw     zero,-44(fp)
'{"PC = 312 : SH", 78, 2740, 16, 32'h7fff0000},         // 00312 sh     a5,-32(fp)
'{"PC = 320 : SB", 80, 2755, 8, 32'h0000000e},          // 00320 sb     a5,-17(fp)
'{"PC = 328 : SB", 82, 2747, 8, 32'h0000000f},          // 00328 sb     a5,-25(fp)
'{"PC = 336 : SB", 84, 2746, 8, 32'h00000001},          // 00336 sb     a5,-26(fp)
'{"PC = 344 : SH", 86, 2744, 16, 32'hfffffffe},         // 00344 sh     a5,-28(fp)
'{"PC = 352 : SH", 88, 2742, 16, 32'h0000000f},         // 00352 sh     a5,-30(fp)
'{"PC = 356 : SH", 89, 2740, 16, 32'h00000000},         // 00356 sh     zero,-32(fp)
'{"PC = 364 : SW", 91, 2736, 32, 32'hfffffffe},         // 00364 sw     a5,-36(fp)
'{"PC = 376 : SW", 94, 2732, 32, 32'h0f0f070f},         // 00376 sw     a5,-40(fp)
'{"PC = 380 : SW", 95, 2728, 32, 32'h00000000},         // 00380 sw     zero,-44(fp)
'{"PC = 396 : SH", 99, 2740, 16, 32'h00000001},         // 00396 sh     a5,-32(fp)
'{"PC = 404 : SB", 101, 2755, 8, 32'h0000000e},         // 00404 sb     a5,-17(fp)
'{"PC = 412 : SB", 103, 2747, 8, 32'h0000000f},         // 00412 sb     a5,-25(fp)
'{"PC = 420 : SB", 105, 2746, 8, 32'h00000001},         // 00420 sb     a5,-26(fp)
'{"PC = 428 : SH", 107, 2744, 16, 32'hfffffffe},                // 00428 sh     a5,-28(fp)
'{"PC = 436 : SH", 109, 2742, 16, 32'h0000000f},                // 00436 sh     a5,-30(fp)
'{"PC = 440 : SH", 110, 2740, 16, 32'h00000000},                // 00440 sh     zero,-32(fp)
'{"PC = 448 : SW", 112, 2736, 32, 32'hfffffffe},                // 00448 sw     a5,-36(fp)
'{"PC = 460 : SW", 115, 2732, 32, 32'h0f0f070f},                // 00460 sw     a5,-40(fp)
'{"PC = 464 : SW", 116, 2728, 32, 32'h00000000},                // 00464 sw     zero,-44(fp)
'{"PC = 480 : SW", 120, 2728, 32, 32'hffffffff},                // 00480 sw     a5,-44(fp)
'{"PC = 488 : SB", 122, 2755, 8, 32'h0000000e},         // 00488 sb     a5,-17(fp)
'{"PC = 496 : SB", 124, 2747, 8, 32'h0000000f},         // 00496 sb     a5,-25(fp)
'{"PC = 504 : SB", 126, 2746, 8, 32'h00000001},         // 00504 sb     a5,-26(fp)
'{"PC = 512 : SH", 128, 2744, 16, 32'hfffffffe},                // 00512 sh     a5,-28(fp)
'{"PC = 520 : SH", 130, 2742, 16, 32'h0000000f},                // 00520 sh     a5,-30(fp)
'{"PC = 524 : SH", 131, 2740, 16, 32'h00000000},                // 00524 sh     zero,-32(fp)
'{"PC = 532 : SW", 133, 2736, 32, 32'hfffffffe},                // 00532 sw     a5,-36(fp)
'{"PC = 544 : SW", 136, 2732, 32, 32'h0f0f070f},                // 00544 sw     a5,-40(fp)
'{"PC = 548 : SW", 137, 2728, 32, 32'h00000000},                // 00548 sw     zero,-44(fp)
'{"PC = 564 : SW", 141, 2728, 32, 32'hf0f0f8f1},                // 00564 sw     a5,-44(fp)
'{"PC = 572 : SB", 143, 2755, 8, 32'h0000000e},         // 00572 sb     a5,-17(fp)
'{"PC = 580 : SB", 145, 2747, 8, 32'h0000000f},         // 00580 sb     a5,-25(fp)
'{"PC = 588 : SB", 147, 2746, 8, 32'h00000001},         // 00588 sb     a5,-26(fp)
'{"PC = 596 : SH", 149, 2744, 16, 32'hfffffffe},                // 00596 sh     a5,-28(fp)
'{"PC = 604 : SH", 151, 2742, 16, 32'h0000000f},                // 00604 sh     a5,-30(fp)
'{"PC = 608 : SH", 152, 2740, 16, 32'h00000000},                // 00608 sh     zero,-32(fp)
'{"PC = 616 : SW", 154, 2736, 32, 32'hfffffffe},                // 00616 sw     a5,-36(fp)
'{"PC = 628 : SW", 157, 2732, 32, 32'h0f0f070f},                // 00628 sw     a5,-40(fp)
'{"PC = 632 : SW", 158, 2728, 32, 32'h00000000},                // 00632 sw     zero,-44(fp)
'{"PC = 652 : SB", 163, 2746, 8, 32'h00000001},         // 00652 sb     a5,-26(fp)
'{"PC = 672 : SH", 168, 2740, 16, 32'h00000000},                // 00672 sh     a5,-32(fp)
'{"PC = 680 : SB", 170, 2755, 8, 32'h0000000e},         // 00680 sb     a5,-17(fp)
'{"PC = 688 : SB", 172, 2747, 8, 32'h0000000f},         // 00688 sb     a5,-25(fp)
'{"PC = 696 : SB", 174, 2746, 8, 32'h00000001},         // 00696 sb     a5,-26(fp)
'{"PC = 704 : SH", 176, 2744, 16, 32'hfffffffe},                // 00704 sh     a5,-28(fp)
'{"PC = 712 : SH", 178, 2742, 16, 32'h0000000f},                // 00712 sh     a5,-30(fp)
'{"PC = 716 : SH", 179, 2740, 16, 32'h00000000},                // 00716 sh     zero,-32(fp)
'{"PC = 724 : SW", 181, 2736, 32, 32'hfffffffe},                // 00724 sw     a5,-36(fp)
'{"PC = 736 : SW", 184, 2732, 32, 32'h0f0f070f},                // 00736 sw     a5,-40(fp)
'{"PC = 740 : SW", 185, 2728, 32, 32'h00000000},                // 00740 sw     zero,-44(fp)
'{"PC = 760 : SB", 190, 2753, 8, 32'h00000001},         // 00760 sb     a5,-19(fp)
'{"PC = 780 : SH", 195, 2746, 16, 32'h00000000},                // 00780 sh     a5,-26(fp)
'{"PC = 788 : SB", 197, 2755, 8, 32'h0000000e},         // 00788 sb     a5,-17(fp)
'{"PC = 796 : SB", 199, 2747, 8, 32'h0000000f},         // 00796 sb     a5,-25(fp)
'{"PC = 804 : SB", 201, 2746, 8, 32'h00000001},         // 00804 sb     a5,-26(fp)
'{"PC = 812 : SH", 203, 2744, 16, 32'hfffffffe},                // 00812 sh     a5,-28(fp)
'{"PC = 820 : SH", 205, 2742, 16, 32'h0000000f},                // 00820 sh     a5,-30(fp)
'{"PC = 824 : SH", 206, 2740, 16, 32'h00000000},                // 00824 sh     zero,-32(fp)
'{"PC = 832 : SW", 208, 2736, 32, 32'hfffffffe},                // 00832 sw     a5,-36(fp)
'{"PC = 844 : SW", 211, 2732, 32, 32'h0f0f070f},                // 00844 sw     a5,-40(fp)
'{"PC = 848 : SW", 212, 2728, 32, 32'h00000000},                // 00848 sw     zero,-44(fp)
'{"PC = 864 : SH", 216, 2740, 16, 32'h00000001},                // 00864 sh     a5,-32(fp)
'{"PC = 872 : SB", 218, 2755, 8, 32'h0000000e},         // 00872 sb     a5,-17(fp)
'{"PC = 880 : SB", 220, 2747, 8, 32'h0000000f},         // 00880 sb     a5,-25(fp)
'{"PC = 888 : SB", 222, 2746, 8, 32'h00000001},         // 00888 sb     a5,-26(fp)
'{"PC = 896 : SH", 224, 2744, 16, 32'hfffffffe},                // 00896 sh     a5,-28(fp)
'{"PC = 904 : SH", 226, 2742, 16, 32'h0000000f},                // 00904 sh     a5,-30(fp)
'{"PC = 908 : SH", 227, 2740, 16, 32'h00000000},                // 00908 sh     zero,-32(fp)
'{"PC = 916 : SW", 229, 2736, 32, 32'hfffffffe},                // 00916 sw     a5,-36(fp)
'{"PC = 928 : SW", 232, 2732, 32, 32'h0f0f070f},                // 00928 sw     a5,-40(fp)
'{"PC = 932 : SW", 233, 2728, 32, 32'h00000000},                // 00932 sw     zero,-44(fp)
'{"PC = 948 : SB", 237, 2746, 8, 32'h00000001},         // 00948 sb     a5,-26(fp)
'{"PC = 964 : SH", 241, 2740, 16, 32'hffff0011},                // 00964 sh     a5,-32(fp)
'{"PC = 972 : SB", 243, 2755, 8, 32'h0000000e},         // 00972 sb     a5,-17(fp)
'{"PC = 980 : SB", 245, 2747, 8, 32'h0000000f},         // 00980 sb     a5,-25(fp)
'{"PC = 988 : SB", 247, 2746, 8, 32'h00000001},         // 00988 sb     a5,-26(fp)
'{"PC = 996 : SH", 249, 2744, 16, 32'hfffffffe},                // 00996 sh     a5,-28(fp)
'{"PC = 1004 : SH", 251, 2742, 16, 32'h0000000f},               // 01004 sh     a5,-30(fp)
'{"PC = 1008 : SH", 252, 2740, 16, 32'h00000000},               // 01008 sh     zero,-32(fp)
'{"PC = 1016 : SW", 254, 2736, 32, 32'hfffffffe},               // 01016 sw     a5,-36(fp)
'{"PC = 1028 : SW", 257, 2732, 32, 32'h0f0f070f},               // 01028 sw     a5,-40(fp)
'{"PC = 1032 : SW", 258, 2728, 32, 32'h00000000},               // 01032 sw     zero,-44(fp)
'{"PC = 1044 : SH", 261, 2740, 16, 32'h001fffc0},               // 01044 sh     a5,-32(fp)
'{"PC = 1056 : SB", 264, 2746, 8, 32'h000001c0},                // 01056 sb     a5,-26(fp)
'{"PC = 1064 : SB", 266, 2755, 8, 32'h0000000e},                // 01064 sb     a5,-17(fp)
'{"PC = 1072 : SB", 268, 2747, 8, 32'h0000000f},                // 01072 sb     a5,-25(fp)
'{"PC = 1080 : SB", 270, 2746, 8, 32'h00000001},                // 01080 sb     a5,-26(fp)
'{"PC = 1088 : SH", 272, 2744, 16, 32'hfffffffe},               // 01088 sh     a5,-28(fp)
'{"PC = 1096 : SH", 274, 2742, 16, 32'h0000000f},               // 01096 sh     a5,-30(fp)
'{"PC = 1100 : SH", 275, 2740, 16, 32'h00000000},               // 01100 sh     zero,-32(fp)
'{"PC = 1108 : SW", 277, 2736, 32, 32'hfffffffe},               // 01108 sw     a5,-36(fp)
'{"PC = 1120 : SW", 280, 2732, 32, 32'h0f0f070f},               // 01120 sw     a5,-40(fp)
'{"PC = 1124 : SW", 281, 2728, 32, 32'h00000000},               // 01124 sw     zero,-44(fp)
'{"PC = 1136 : SH", 284, 2755, 16, 32'h00007f87},               // 01136 sh     a5,-17(fp)
'{"PC = 1148 : SB", 287, 2746, 8, 32'h00000010},                // 01148 sb     a5,-26(fp)
'{"PC = 1156 : SB", 289, 2755, 8, 32'h0000000e},                // 01156 sb     a5,-17(fp)
'{"PC = 1164 : SB", 291, 2747, 8, 32'h0000000f},                // 01164 sb     a5,-25(fp)
'{"PC = 1172 : SB", 293, 2746, 8, 32'h00000001},                // 01172 sb     a5,-26(fp)
'{"PC = 1180 : SH", 295, 2744, 16, 32'hfffffffe},               // 01180 sh     a5,-28(fp)
'{"PC = 1188 : SH", 297, 2742, 16, 32'h0000000f},               // 01188 sh     a5,-30(fp)
'{"PC = 1192 : SH", 298, 2740, 16, 32'h00000000},               // 01192 sh     zero,-32(fp)
'{"PC = 1200 : SW", 300, 2736, 32, 32'hfffffffe},               // 01200 sw     a5,-36(fp)
'{"PC = 1212 : SW", 303, 2732, 32, 32'h0f0f070f},               // 01212 sw     a5,-40(fp)
'{"PC = 1216 : SW", 304, 2728, 32, 32'h00000000},               // 01216 sw     zero,-44(fp)
'{"PC = 1236 : SW", 309, 2728, 32, 32'h0000070f},               // 01236 sw     a4,-44(fp)
'{"PC = 1240 : SW", 310, 2732, 32, 32'h000007ff},               // 01240 sw     a5,-40(fp)
'{"PC = 1248 : SB", 312, 2755, 8, 32'h0000000e},                // 01248 sb     a5,-17(fp)
'{"PC = 1256 : SB", 314, 2747, 8, 32'h0000000f},                // 01256 sb     a5,-25(fp)
'{"PC = 1264 : SB", 316, 2746, 8, 32'h00000001},                // 01264 sb     a5,-26(fp)
'{"PC = 1272 : SH", 318, 2744, 16, 32'hfffffffe},               // 01272 sh     a5,-28(fp)
'{"PC = 1280 : SH", 320, 2742, 16, 32'h0000000f},               // 01280 sh     a5,-30(fp)
'{"PC = 1284 : SH", 321, 2740, 16, 32'h00000000},               // 01284 sh     zero,-32(fp)
'{"PC = 1292 : SW", 323, 2736, 32, 32'hfffffffe},               // 01292 sw     a5,-36(fp)
'{"PC = 1304 : SW", 326, 2732, 32, 32'h0f0f070f},               // 01304 sw     a5,-40(fp)
'{"PC = 1308 : SW", 327, 2728, 32, 32'h00000000},               // 01308 sw     zero,-44(fp)
'{"PC = 1328 : SW", 332, 2728, 32, 32'hf0f0f8f1},               // 01328 sw     a5,-44(fp)
'{"PC = 1348 : SB", 337, 2755, 8, 32'h0000000e},                // 01348 sb     a5,-17(fp)
'{"PC = 1356 : SB", 339, 2747, 8, 32'h0000000f},                // 01356 sb     a5,-25(fp)
'{"PC = 1364 : SB", 341, 2746, 8, 32'h00000001},                // 01364 sb     a5,-26(fp)
'{"PC = 1372 : SH", 343, 2744, 16, 32'hfffffffe},               // 01372 sh     a5,-28(fp)
'{"PC = 1380 : SH", 345, 2742, 16, 32'h0000000f},               // 01380 sh     a5,-30(fp)
'{"PC = 1384 : SH", 346, 2740, 16, 32'h00000000},               // 01384 sh     zero,-32(fp)
'{"PC = 1392 : SW", 348, 2736, 32, 32'hfffffffe},               // 01392 sw     a5,-36(fp)
'{"PC = 1404 : SW", 351, 2732, 32, 32'h0f0f070f},               // 01404 sw     a5,-40(fp)
'{"PC = 1408 : SW", 352, 2728, 32, 32'h00000000},               // 01408 sw     zero,-44(fp)
'{"PC = 1424 : SB", 356, 2746, 8, 32'h00000001},                // 01424 sb     a5,-26(fp)
'{"PC = 1440 : SH", 360, 2740, 16, 32'h00000000},               // 01440 sh     a5,-32(fp)
'{"PC = 1448 : SB", 362, 2755, 8, 32'h0000000e},                // 01448 sb     a5,-17(fp)
'{"PC = 1456 : SB", 364, 2747, 8, 32'h0000000f},                // 01456 sb     a5,-25(fp)
'{"PC = 1464 : SB", 366, 2746, 8, 32'h00000001},                // 01464 sb     a5,-26(fp)
'{"PC = 1472 : SH", 368, 2744, 16, 32'hfffffffe},               // 01472 sh     a5,-28(fp)
'{"PC = 1480 : SH", 370, 2742, 16, 32'h0000000f},               // 01480 sh     a5,-30(fp)
'{"PC = 1484 : SH", 371, 2740, 16, 32'h00000000},               // 01484 sh     zero,-32(fp)
'{"PC = 1492 : SW", 373, 2736, 32, 32'hfffffffe},               // 01492 sw     a5,-36(fp)
'{"PC = 1504 : SW", 376, 2732, 32, 32'h0f0f070f},               // 01504 sw     a5,-40(fp)
'{"PC = 1508 : SW", 377, 2728, 32, 32'h00000000},               // 01508 sw     zero,-44(fp)
'{"PC = 1524 : SH", 381, 2746, 16, 32'h00000001},               // 01524 sh     a5,-26(fp)
'{"PC = 1540 : SH", 385, 2740, 16, 32'h00000000},               // 01540 sh     a5,-32(fp)
'{"PC = 1548 : SB", 387, 2755, 8, 32'h0000000e},                // 01548 sb     a5,-17(fp)
'{"PC = 1556 : SB", 389, 2747, 8, 32'h0000000f},                // 01556 sb     a5,-25(fp)
'{"PC = 1564 : SB", 391, 2746, 8, 32'h00000001},                // 01564 sb     a5,-26(fp)
'{"PC = 1572 : SH", 393, 2744, 16, 32'hfffffffe},               // 01572 sh     a5,-28(fp)
'{"PC = 1580 : SH", 395, 2742, 16, 32'h0000000f},               // 01580 sh     a5,-30(fp)
'{"PC = 1584 : SH", 396, 2740, 16, 32'h00000000},               // 01584 sh     zero,-32(fp)
'{"PC = 1592 : SW", 398, 2736, 32, 32'hfffffffe},               // 01592 sw     a5,-36(fp)
'{"PC = 1604 : SW", 401, 2732, 32, 32'h0f0f070f},               // 01604 sw     a5,-40(fp)
'{"PC = 1608 : SW", 402, 2728, 32, 32'h00000000},               // 01608 sw     zero,-44(fp)
'{"PC = 1620 : SH", 405, 2740, 16, 32'h00000001},               // 01620 sh     a5,-32(fp)
'{"PC = 1628 : SB", 407, 2755, 8, 32'h0000000e},                // 01628 sb     a5,-17(fp)
'{"PC = 1636 : SB", 409, 2747, 8, 32'h0000000f},                // 01636 sb     a5,-25(fp)
'{"PC = 1644 : SB", 411, 2746, 8, 32'h00000001},                // 01644 sb     a5,-26(fp)
'{"PC = 1652 : SH", 413, 2744, 16, 32'hfffffffe},               // 01652 sh     a5,-28(fp)
'{"PC = 1660 : SH", 415, 2742, 16, 32'h0000000f},               // 01660 sh     a5,-30(fp)
'{"PC = 1664 : SH", 416, 2740, 16, 32'h00000000},               // 01664 sh     zero,-32(fp)
'{"PC = 1672 : SW", 418, 2736, 32, 32'hfffffffe},               // 01672 sw     a5,-36(fp)
'{"PC = 1684 : SW", 421, 2732, 32, 32'h0f0f070f},               // 01684 sw     a5,-40(fp)
'{"PC = 1688 : SW", 422, 2728, 32, 32'h00000000},               // 01688 sw     zero,-44(fp)
'{"PC = 1724 : SB", 430, 2755, 8, 32'h0000000e},                // 01724 sb     a5,-17(fp)
'{"PC = 1732 : SB", 432, 2755, 8, 32'h0000000e},                // 01732 sb     a5,-17(fp)
'{"PC = 1740 : SB", 434, 2747, 8, 32'h0000000f},                // 01740 sb     a5,-25(fp)
'{"PC = 1748 : SB", 436, 2746, 8, 32'h00000001},                // 01748 sb     a5,-26(fp)
'{"PC = 1756 : SH", 438, 2744, 16, 32'hfffffffe},               // 01756 sh     a5,-28(fp)
'{"PC = 1764 : SH", 440, 2742, 16, 32'h0000000f},               // 01764 sh     a5,-30(fp)
'{"PC = 1768 : SH", 441, 2740, 16, 32'h00000000},               // 01768 sh     zero,-32(fp)
'{"PC = 1776 : SW", 443, 2736, 32, 32'hfffffffe},               // 01776 sw     a5,-36(fp)
'{"PC = 1788 : SW", 446, 2732, 32, 32'h0f0f070f},               // 01788 sw     a5,-40(fp)
'{"PC = 1792 : SW", 447, 2728, 32, 32'h00000000},               // 01792 sw     zero,-44(fp)
'{"PC = 1828 : SB", 456, 2755, 8, 32'h00000000},                // 01828 sb     a5,-17(fp)
'{"PC = 1836 : SB", 458, 2755, 8, 32'h0000000e},                // 01836 sb     a5,-17(fp)
'{"PC = 1844 : SB", 460, 2747, 8, 32'h0000000f},                // 01844 sb     a5,-25(fp)
'{"PC = 1852 : SB", 462, 2746, 8, 32'h00000001},                // 01852 sb     a5,-26(fp)
'{"PC = 1860 : SH", 464, 2744, 16, 32'hfffffffe},               // 01860 sh     a5,-28(fp)
'{"PC = 1868 : SH", 466, 2742, 16, 32'h0000000f},               // 01868 sh     a5,-30(fp)
'{"PC = 1872 : SH", 467, 2740, 16, 32'h00000000},               // 01872 sh     zero,-32(fp)
'{"PC = 1880 : SW", 469, 2736, 32, 32'hfffffffe},               // 01880 sw     a5,-36(fp)
'{"PC = 1892 : SW", 472, 2732, 32, 32'h0f0f070f},               // 01892 sw     a5,-40(fp)
'{"PC = 1896 : SW", 473, 2728, 32, 32'h00000000},               // 01896 sw     zero,-44(fp)
'{"PC = 1928 : SB", 481, 2755, 8, 32'h00000000},                // 01928 sb     zero,-17(fp)
'{"PC = 1936 : SB", 483, 2755, 8, 32'h0000000e},                // 01936 sb     a5,-17(fp)
'{"PC = 1944 : SB", 485, 2747, 8, 32'h0000000f},                // 01944 sb     a5,-25(fp)
'{"PC = 1952 : SB", 487, 2746, 8, 32'h00000001},                // 01952 sb     a5,-26(fp)
'{"PC = 1960 : SH", 489, 2744, 16, 32'hfffffffe},               // 01960 sh     a5,-28(fp)
'{"PC = 1968 : SH", 491, 2742, 16, 32'h0000000f},               // 01968 sh     a5,-30(fp)
'{"PC = 1972 : SH", 492, 2740, 16, 32'h00000000},               // 01972 sh     zero,-32(fp)
'{"PC = 1980 : SW", 494, 2736, 32, 32'hfffffffe},               // 01980 sw     a5,-36(fp)
'{"PC = 1992 : SW", 497, 2732, 32, 32'h0f0f070f},               // 01992 sw     a5,-40(fp)
'{"PC = 1996 : SW", 498, 2728, 32, 32'h00000000},               // 01996 sw     zero,-44(fp)
'{"PC = 2028 : SB", 506, 2755, 8, 32'h00000000},                // 02028 sb     zero,-17(fp)
'{"PC = 2036 : SB", 508, 2755, 8, 32'h0000000e},                // 02036 sb     a5,-17(fp)
'{"PC = 2044 : SB", 510, 2747, 8, 32'h0000000f},                // 02044 sb     a5,-25(fp)
'{"PC = 2052 : SB", 512, 2746, 8, 32'h00000001},                // 02052 sb     a5,-26(fp)
'{"PC = 2060 : SH", 514, 2744, 16, 32'hfffffffe},               // 02060 sh     a5,-28(fp)
'{"PC = 2068 : SH", 516, 2742, 16, 32'h0000000f},               // 02068 sh     a5,-30(fp)
'{"PC = 2072 : SH", 517, 2740, 16, 32'h00000000},               // 02072 sh     zero,-32(fp)
'{"PC = 2080 : SW", 519, 2736, 32, 32'hfffffffe},               // 02080 sw     a5,-36(fp)
'{"PC = 2092 : SW", 522, 2732, 32, 32'h0f0f070f},               // 02092 sw     a5,-40(fp)
'{"PC = 2096 : SW", 523, 2728, 32, 32'h00000000},               // 02096 sw     zero,-44(fp)
'{"PC = 2128 : SB", 531, 2755, 8, 32'h00000000},                // 02128 sb     zero,-17(fp)
'{"PC = 2136 : SB", 533, 2755, 8, 32'h0000000e},                // 02136 sb     a5,-17(fp)
'{"PC = 2144 : SB", 535, 2747, 8, 32'h0000000f},                // 02144 sb     a5,-25(fp)
'{"PC = 2152 : SB", 537, 2746, 8, 32'h00000001},                // 02152 sb     a5,-26(fp)
'{"PC = 2160 : SH", 539, 2744, 16, 32'hfffffffe},               // 02160 sh     a5,-28(fp)
'{"PC = 2168 : SH", 541, 2742, 16, 32'h0000000f},               // 02168 sh     a5,-30(fp)
'{"PC = 2172 : SH", 542, 2740, 16, 32'h00000000},               // 02172 sh     zero,-32(fp)
'{"PC = 2180 : SW", 544, 2736, 32, 32'hfffffffe},               // 02180 sw     a5,-36(fp)
'{"PC = 2192 : SW", 547, 2732, 32, 32'h0f0f070f},               // 02192 sw     a5,-40(fp)
'{"PC = 2196 : SW", 548, 2728, 32, 32'h00000000},               // 02196 sw     zero,-44(fp)
'{"PC = 2228 : SB", 556, 2755, 8, 32'h00000000},                // 02228 sb     zero,-17(fp)
'{"PC = 2236 : SB", 558, 2755, 8, 32'h0000000e},                // 02236 sb     a5,-17(fp)
'{"PC = 2244 : SB", 560, 2747, 8, 32'h0000000f},                // 02244 sb     a5,-25(fp)
'{"PC = 2252 : SB", 562, 2746, 8, 32'h00000001},                // 02252 sb     a5,-26(fp)
'{"PC = 2260 : SH", 564, 2744, 16, 32'hfffffffe},               // 02260 sh     a5,-28(fp)
'{"PC = 2268 : SH", 566, 2742, 16, 32'h0000000f},               // 02268 sh     a5,-30(fp)
'{"PC = 2272 : SH", 567, 2740, 16, 32'h00000000},               // 02272 sh     zero,-32(fp)
'{"PC = 2280 : SW", 569, 2736, 32, 32'hfffffffe},               // 02280 sw     a5,-36(fp)
'{"PC = 2292 : SW", 572, 2732, 32, 32'h0f0f070f},               // 02292 sw     a5,-40(fp)
'{"PC = 2296 : SW", 573, 2728, 32, 32'h00000000},               // 02296 sw     zero,-44(fp)
'{"PC = 2308 : SW", 576, 2732, 32, 32'h00000000},               // 02308 sw     a4,-40(fp)
'{"PC = 2316 : SB", 578, 2755, 8, 32'h0000000e},                // 02316 sb     a5,-17(fp)
'{"PC = 2324 : SB", 580, 2747, 8, 32'h0000000f},                // 02324 sb     a5,-25(fp)
'{"PC = 2332 : SB", 582, 2746, 8, 32'h00000001},                // 02332 sb     a5,-26(fp)
'{"PC = 2340 : SH", 584, 2744, 16, 32'hfffffffe},               // 02340 sh     a5,-28(fp)
'{"PC = 2348 : SH", 586, 2742, 16, 32'h0000000f},               // 02348 sh     a5,-30(fp)
'{"PC = 2352 : SH", 587, 2740, 16, 32'h00000000},               // 02352 sh     zero,-32(fp)
'{"PC = 2360 : SW", 589, 2736, 32, 32'hfffffffe},               // 02360 sw     a5,-36(fp)
'{"PC = 2372 : SW", 592, 2732, 32, 32'h0f0f070f},               // 02372 sw     a5,-40(fp)
'{"PC = 2376 : SW", 593, 2728, 32, 32'h00000000},               // 02376 sw     zero,-44(fp)
'{"PC = 2388 : SW", 596, 2732, 32, 32'h0000e950},               // 02388 sw     a4,-40(fp)
'{"PC = 2396 : SB", 598, 2755, 8, 32'h0000000e},                // 02396 sb     a5,-17(fp)
'{"PC = 2404 : SB", 600, 2747, 8, 32'h0000000f},                // 02404 sb     a5,-25(fp)
'{"PC = 2412 : SB", 602, 2746, 8, 32'h00000001},                // 02412 sb     a5,-26(fp)
'{"PC = 2420 : SH", 604, 2744, 16, 32'hfffffffe},               // 02420 sh     a5,-28(fp)
'{"PC = 2428 : SH", 606, 2742, 16, 32'h0000000f},               // 02428 sh     a5,-30(fp)
'{"PC = 2432 : SH", 607, 2740, 16, 32'h00000000},               // 02432 sh     zero,-32(fp)
'{"PC = 2440 : SW", 609, 2736, 32, 32'hfffffffe},               // 02440 sw     a5,-36(fp)
'{"PC = 2452 : SW", 612, 2732, 32, 32'h0f0f070f},               // 02452 sw     a5,-40(fp)
'{"PC = 2456 : SW", 613, 2728, 32, 32'h00000000},               // 02456 sw     zero,-44(fp)
'{"PC = 2460 : SB", 614, 2755, 8, 32'h00000000},                // 02460 sb     zero,-17(fp)
'{"PC = 2464 : SW", 615, 2748, 32, 32'h00000000},               // 02464 sw     zero,-24(fp)
'{"PC = 2496 : SB", 630, 2755, 8, 32'h00000001},                // 02496 sb     a5,-17(fp)
'{"PC = 2508 : SW", 633, 2748, 32, 32'h00000001},               // 02508 sw     a5,-24(fp)
'{"PC = 2540 : SW", 641, 2732, 32, 32'h00000000},               // 02540 sw     t1,-40(fp)
'{"PC = 2548 : SB", 643, 2755, 8, 32'h0000000e},                // 02548 sb     a5,-17(fp)
'{"PC = 2556 : SB", 645, 2747, 8, 32'h0000000f},                // 02556 sb     a5,-25(fp)
'{"PC = 2564 : SB", 647, 2746, 8, 32'h00000001},                // 02564 sb     a5,-26(fp)
'{"PC = 2572 : SH", 649, 2744, 16, 32'hfffffffe},               // 02572 sh     a5,-28(fp)
'{"PC = 2580 : SH", 651, 2742, 16, 32'h0000000f},               // 02580 sh     a5,-30(fp)
'{"PC = 2584 : SH", 652, 2740, 16, 32'h00000000},               // 02584 sh     zero,-32(fp)
'{"PC = 2592 : SW", 654, 2736, 32, 32'hfffffffe},               // 02592 sw     a5,-36(fp)
'{"PC = 2604 : SW", 657, 2732, 32, 32'h0f0f070f},               // 02604 sw     a5,-40(fp)
'{"PC = 2608 : SW", 658, 2728, 32, 32'h00000000},               // 02608 sw     zero,-44(fp)
'{"PC = 2644 : SB", 666, 2755, 8, 32'h0000000e},                // 02644 sb     a5,-17(fp)
'{"PC = 2652 : SB", 668, 2747, 8, 32'h0000000f},                // 02652 sb     a5,-25(fp)
'{"PC = 2660 : SB", 670, 2746, 8, 32'h00000001},                // 02660 sb     a5,-26(fp)
'{"PC = 2668 : SH", 672, 2744, 16, 32'hfffffffe},               // 02668 sh     a5,-28(fp)
'{"PC = 2676 : SH", 674, 2742, 16, 32'h0000000f},               // 02676 sh     a5,-30(fp)
'{"PC = 2680 : SH", 675, 2740, 16, 32'h00000000},               // 02680 sh     zero,-32(fp)
'{"PC = 2688 : SW", 677, 2736, 32, 32'hfffffffe},               // 02688 sw     a5,-36(fp)
'{"PC = 2700 : SW", 680, 2732, 32, 32'h0f0f070f},               // 02700 sw     a5,-40(fp)
'{"PC = 2704 : SW", 681, 2728, 32, 32'h00000000}                // 02704 sw     zero,-44(fp)
};

bit clk;
bit reset;

// Design Under Test
riscv #(MEM_SIZE) riscv1 (
    .clk(clk),
    .rst(reset)
);

initial $timeformat ( -9, 1, " ns", 12 );

// Clock and Reset Definitin
initial begin
    clk = 1'b1;
    reset = 1'b1;
    #(CLK_PERIOD) reset = 1'b0;
end

always
    #(CLK_PERIOD/2) clk = ~clk;

// Load the program in the instruction memory from a binary file
initial begin
    // Init the memory with 0
    for (int i = 0; i < MEM_SIZE+1; i=i+1) begin
        riscv1.mem1.mem[i] = 8'hff;
    end
    $readmemb("D:/Dossier principal/Electronique/Tout MES programmes/RISC_V_Project/prog/asm_bench_global.bin", insn_buff);
    for (int i = 0; i < PROG_SIZE; i=i+1) begin
        riscv1.mem1.mem[4*i  ] = insn_buff[i][7:0];
        riscv1.mem1.mem[4*i+1] = insn_buff[i][15:8];
        riscv1.mem1.mem[4*i+2] = insn_buff[i][23:16];
        riscv1.mem1.mem[4*i+3] = insn_buff[i][31:24];
    end
    
    clk <= 1'b0  ;
    reset <= 1'b1;
    #21 reset <= 1'b0;
    clock_number = 0;
end

always @(posedge clk) begin
    clock_number = clock_number + 1;
    
    //----- Tests généraux
    for (int i = 0; i < NB_TESTS; i++) begin
        if (clock_number == test[i].clk+5) begin      // +5 because of the stages of the pipeline
        // if (clock_number == test[i].clk+4) begin      // +4 because of the stages of the pipeline
            $display("========== Test %s (CLK = %d)", test[i].name, clock_number);
            $display("Expected value : 0x%h @ 0x%h",  test[i].value, test[i].address);
            value_ok = 0;
            case (test[i].size)
                8: begin
                    $display(
                        "Read value     : 0x%h @ 0x%h", 
                        riscv1.mem1.mem[test[i].address], 
                        test[i].address
                    );
                    if (riscv1.mem1.mem[test[i].address  ][7:0]  == test[i].value[7:0]) begin
                        value_ok = 1;
                    end
                end
                16: begin
                    $display(
                        "Read value     : 0x%h %h @ 0x%h", 
                        riscv1.mem1.mem[test[i].address+1], 
                        riscv1.mem1.mem[test[i].address], 
                        test[i].address
                    );
                    if (riscv1.mem1.mem[test[i].address  ][7:0]  == test[i].value[7:0] &&
                        riscv1.mem1.mem[test[i].address+1][7:0]  == test[i].value[15:8]) begin
                        value_ok = 1;
                    end
                end
                32: begin
                    $display(
                        "Read value     : 0x%h %h %h %h @ 0x%h", 
                        riscv1.mem1.mem[test[i].address+3], 
                        riscv1.mem1.mem[test[i].address+2], 
                        riscv1.mem1.mem[test[i].address+1], 
                        riscv1.mem1.mem[test[i].address], 
                        test[i].address
                    );
                    if (riscv1.mem1.mem[test[i].address  ][7:0]  == test[i].value[7:0] &&
                        riscv1.mem1.mem[test[i].address+1][7:0]  == test[i].value[15:8] &&
                        riscv1.mem1.mem[test[i].address+2][7:0]  == test[i].value[23:16] &&
                        riscv1.mem1.mem[test[i].address+3][7:0]  == test[i].value[31:24]) begin
                        value_ok = 1;
                    end
                end
                default: begin
                    $display("ERROR : Wrong size");
                    $finish;
                end
            endcase
            if (value_ok == 0) begin
                $display("ERROR : Expected value is not the same as the read value");
                // $finish;
            end
            else begin
                $display("TEST PASSED");
                passed_test = passed_test + 1;
            end
            done_test = done_test + 1;
        end
    end
    if (done_test == NB_TESTS) begin
        $display("");
        $display("========== %d tests passed on %d", passed_test, done_test);
        // $finish;
    end
end
endmodule